module Comparator_tb;
reg [31:0] a;
reg [31:0] b;
reg [2:0] op;

wire compout;

//op=000 a==b
//op=001 a>=b
//op=010 a<=b
//op=011 a>b
//op=100 a<b
//op=101 a!=b

Comparator dut (a, b, op, compout);
initial
	begin
	$dumpfile("saidaComparator.vcd"); //Serve para olhar pelo gtkwave, sinal de onda. Basta dar: gtkwave saidaComparator.vcd
	$dumpvars;
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b000;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b000;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b001;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b001;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000001;
	b = 32'b00000000000000000000000000000000;
	op= 3'b001;
	$display(compout);
	#10
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b010;
	$display(compout);
	#10
	a = 32'b00000000000000000000000000000001;
	b = 32'b00000000000000000000000000000000;
	op= 3'b010;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b010;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b011;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000001;
	b = 32'b00000000000000000000000000000000;
	op= 3'b011;
	$display(compout);
	#10
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b011;
	$display(compout);
	#10
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b100;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000001;
	b = 32'b00000000000000000000000000000000;
	op= 3'b100;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b100;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000000;
	op= 3'b101;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000001;
	b = 32'b00000000000000000000000000000000;
	op= 3'b101;
	#10
	$display(compout);
	a = 32'b00000000000000000000000000000000;
	b = 32'b00000000000000000000000000000001;
	op= 3'b101;
	#10
	$display(compout);
	$finish;
	end
endmodule
